library ieee;
use ieee.std_logic_1164.all;

entity divCounter is
	
	port (
	clr: in std_logic;
	clk: in std_logic;
	rxf: out std_logic
	);

end divCounter;
	


